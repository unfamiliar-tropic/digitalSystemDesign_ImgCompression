`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2017/12/18 16:28:02
// Design Name: 
// Module Name: memory_model
// Project Name: 
// Target Devices: 
// Tool Versionext_state: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////




module memory_model(clk, rst, start, finish_ack, data_out, finish, data_all_out, data_start, index1, index2);

    parameter N = 16;
    parameter W = 8;
    
    //number of data line
    parameter D = 4;
	 parameter LOGD = 3;
	
    parameter WAIT = 50;
    parameter LOGWAIT = 7;
    input clk, rst;
	 input start;
    input finish_ack;
    
    output [N*W-1:0] data_out;
    output reg finish;
    output reg data_all_out;
	 output reg data_start;
	 
	 output index1, index2;
    
    //memory 
    reg [W-1:0] data[D-1:0][N-1:0];
    reg[LOGD:0] index;
    reg[LOGWAIT:0] count;
	 
	 assign indexi = index[0];
	 assign index2 = index[1];
    
    reg [1:0] present_state, next_state;
    parameter idle = 2'b00, waiting = 2'b01, data_ready = 2'b10, done = 2'b11;
    
    assign data_out
    	= {data[index][0],data[index][1],data[index][2],data[index][3],data[index][4],data[index][5],data[index][6],data[index][7], 
    		data[index][8],data[index][9],data[index][10],data[index][11],data[index][12],data[index][13],data[index][14],data[index][15]};
    		
    always @(posedge clk or negedge rst) 
        if (!rst) present_state <= idle;
        else present_state <= next_state;
    
    always @(*) case(present_state)

    	idle : 
    		if(start) next_state = waiting;
    		else next_state = idle;
    	
    	waiting :
    		if(count == 0) next_state = data_ready;
    		else next_state = waiting;
    	
    	data_ready :
    		if(finish_ack) begin
				if(index == D-1) next_state = done;
				else next_state = waiting;
			end
		
		done : next_state = done;
    
    endcase
    
    always @(posedge clk or negedge rst) begin
		
		if(!rst) begin
			finish <= 0;
			index <= 0;
			data_all_out <= 0;
			data_start <= 0;
		end
		
		else case(present_state)
			idle : 
				if(start) begin
					finish <= 0;
					count <= WAIT;
					data_all_out <= 0;
					data_start <= 1;
				end
			
			waiting :
				if(count != 0) count <= count-1;
				else begin
					finish <= 1;
				end
			
			data_ready :
				if(finish_ack) begin
					if(index == D-1) begin
						data_all_out <= 1;
						finish <= 0;
					end
					else begin
						finish <= 0;
						index <= index + 1;
						count <= WAIT;
					end
				end
			
			done : ;
				
		endcase
    end
    
    
    
    always @(negedge rst) begin
        /*
    data[0][0] <=10;	data[1][0] <=38;	data[2][0] <=209;	data[3][0] <=9;	data[4][0] <=170;	data[5][0] <=63;	data[6][0] <=228;	data[7][0] <=43;	data[8][0] <=33;	data[9][0] <=113;	data[10][0] <=198;	data[11][0] <=25;	data[12][0] <=233;	data[13][0] <=68;	data[14][0] <=213;	data[15][0] <=246;	data[16][0] <=220;	data[17][0] <=142;	data[18][0] <=91;	data[19][0] <=174;	data[20][0] <=154;	data[21][0] <=199;	data[22][0] <=131;	data[23][0] <=206;	data[24][0] <=12;	data[25][0] <=167;	data[26][0] <=158;	data[27][0] <=3;	data[28][0] <=39;	data[29][0] <=30;	data[30][0] <=74;	data[31][0] <=229;
    data[0][1] <=129;	data[1][1] <=38;	data[2][1] <=211;	data[3][1] <=19;	data[4][1] <=214;	data[5][1] <=231;	data[6][1] <=141;	data[7][1] <=152;	data[8][1] <=40;	data[9][1] <=29;	data[10][1] <=180;	data[11][1] <=58;	data[12][1] <=116;	data[13][1] <=112;	data[14][1] <=244;	data[15][1] <=197;	data[16][1] <=217;	data[17][1] <=53;	data[18][1] <=57;	data[19][1] <=107;	data[20][1] <=84;	data[21][1] <=127;	data[22][1] <=144;	data[23][1] <=216;	data[24][1] <=47;	data[25][1] <=221;	data[26][1] <=124;	data[27][1] <=54;	data[28][1] <=88;	data[29][1] <=15;	data[30][1] <=180;	data[31][1] <=148;
    data[0][2] <=95;	data[1][2] <=2;	data[2][2] <=200;	data[3][2] <=218;	data[4][2] <=40;	data[5][2] <=72;	data[6][2] <=181;	data[7][2] <=172;	data[8][2] <=99;	data[9][2] <=150;	data[10][2] <=206;	data[11][2] <=141;	data[12][2] <=6;	data[13][2] <=183;	data[14][2] <=65;	data[15][2] <=246;	data[16][2] <=11;	data[17][2] <=59;	data[18][2] <=172;	data[19][2] <=204;	data[20][2] <=14;	data[21][2] <=11;	data[22][2] <=204;	data[23][2] <=7;	data[24][2] <=65;	data[25][2] <=204;	data[26][2] <=168;	data[27][2] <=105;	data[28][2] <=47;	data[29][2] <=42;	data[30][2] <=147;	data[31][2] <=246;
    data[0][3] <=65;	data[1][3] <=18;	data[2][3] <=11;	data[3][3] <=52;	data[4][3] <=77;	data[5][3] <=91;	data[6][3] <=227;	data[7][3] <=205;	data[8][3] <=140;	data[9][3] <=235;	data[10][3] <=178;	data[11][3] <=177;	data[12][3] <=128;	data[13][3] <=49;	data[14][3] <=127;	data[15][3] <=183;	data[16][3] <=64;	data[17][3] <=74;	data[18][3] <=173;	data[19][3] <=105;	data[20][3] <=2;	data[21][3] <=36;	data[22][3] <=143;	data[23][3] <=25;	data[24][3] <=150;	data[25][3] <=245;	data[26][3] <=28;	data[27][3] <=116;	data[28][3] <=113;	data[29][3] <=143;	data[30][3] <=154;	data[31][3] <=56;
    data[0][4] <=179;	data[1][4] <=207;	data[2][4] <=54;	data[3][4] <=252;	data[4][4] <=43;	data[5][4] <=155;	data[6][4] <=114;	data[7][4] <=78;	data[8][4] <=17;	data[9][4] <=39;	data[10][4] <=110;	data[11][4] <=138;	data[12][4] <=151;	data[13][4] <=54;	data[14][4] <=159;	data[15][4] <=149;	data[16][4] <=190;	data[17][4] <=231;	data[18][4] <=117;	data[19][4] <=129;	data[20][4] <=38;	data[21][4] <=131;	data[22][4] <=29;	data[23][4] <=83;	data[24][4] <=32;	data[25][4] <=51;	data[26][4] <=182;	data[27][4] <=215;	data[28][4] <=224;	data[29][4] <=222;	data[30][4] <=69;	data[31][4] <=159;
    data[0][5] <=209;	data[1][5] <=74;	data[2][5] <=200;	data[3][5] <=13;	data[4][5] <=65;	data[5][5] <=237;	data[6][5] <=68;	data[7][5] <=150;	data[8][5] <=179;	data[9][5] <=132;	data[10][5] <=151;	data[11][5] <=115;	data[12][5] <=76;	data[13][5] <=51;	data[14][5] <=46;	data[15][5] <=79;	data[16][5] <=123;	data[17][5] <=122;	data[18][5] <=27;	data[19][5] <=121;	data[20][5] <=211;	data[21][5] <=183;	data[22][5] <=8;	data[23][5] <=116;	data[24][5] <=249;	data[25][5] <=171;	data[26][5] <=225;	data[27][5] <=172;	data[28][5] <=79;	data[29][5] <=41;	data[30][5] <=23;	data[31][5] <=233;
    data[0][6] <=108;	data[1][6] <=167;	data[2][6] <=2;	data[3][6] <=32;	data[4][6] <=151;	data[5][6] <=239;	data[6][6] <=59;	data[7][6] <=55;	data[8][6] <=37;	data[9][6] <=45;	data[10][6] <=234;	data[11][6] <=91;	data[12][6] <=227;	data[13][6] <=204;	data[14][6] <=187;	data[15][6] <=224;	data[16][6] <=37;	data[17][6] <=125;	data[18][6] <=109;	data[19][6] <=52;	data[20][6] <=92;	data[21][6] <=109;	data[22][6] <=39;	data[23][6] <=75;	data[24][6] <=26;	data[25][6] <=220;	data[26][6] <=62;	data[27][6] <=22;	data[28][6] <=60;	data[29][6] <=106;	data[30][6] <=37;	data[31][6] <=156;
    data[0][7] <=76;	data[1][7] <=41;	data[2][7] <=84;	data[3][7] <=128;	data[4][7] <=133;	data[5][7] <=194;	data[6][7] <=73;	data[7][7] <=167;	data[8][7] <=152;	data[9][7] <=159;	data[10][7] <=24;	data[11][7] <=94;	data[12][7] <=168;	data[13][7] <=234;	data[14][7] <=147;	data[15][7] <=112;	data[16][7] <=25;	data[17][7] <=55;	data[18][7] <=227;	data[19][7] <=76;	data[20][7] <=94;	data[21][7] <=112;	data[22][7] <=193;	data[23][7] <=119;	data[24][7] <=25;	data[25][7] <=64;	data[26][7] <=163;	data[27][7] <=229;	data[28][7] <=73;	data[29][7] <=203;	data[30][7] <=155;	data[31][7] <=192;
    data[0][8] <=93;	data[1][8] <=42;	data[2][8] <=31;	data[3][8] <=137;	data[4][8] <=82;	data[5][8] <=134;	data[6][8] <=170;	data[7][8] <=143;	data[8][8] <=117;	data[9][8] <=33;	data[10][8] <=228;	data[11][8] <=159;	data[12][8] <=27;	data[13][8] <=182;	data[14][8] <=242;	data[15][8] <=169;	data[16][8] <=35;	data[17][8] <=172;	data[18][8] <=57;	data[19][8] <=204;	data[20][8] <=127;	data[21][8] <=3;	data[22][8] <=205;	data[23][8] <=86;	data[24][8] <=233;	data[25][8] <=101;	data[26][8] <=37;	data[27][8] <=72;	data[28][8] <=172;	data[29][8] <=79;	data[30][8] <=202;	data[31][8] <=33;
    data[0][9] <=206;	data[1][9] <=180;	data[2][9] <=218;	data[3][9] <=31;	data[4][9] <=189;	data[5][9] <=27;	data[6][9] <=71;	data[7][9] <=70;	data[8][9] <=68;	data[9][9] <=242;	data[10][9] <=217;	data[11][9] <=96;	data[12][9] <=172;	data[13][9] <=216;	data[14][9] <=22;	data[15][9] <=156;	data[16][9] <=212;	data[17][9] <=210;	data[18][9] <=45;	data[19][9] <=113;	data[20][9] <=244;	data[21][9] <=163;	data[22][9] <=180;	data[23][9] <=46;	data[24][9] <=237;	data[25][9] <=64;	data[26][9] <=192;	data[27][9] <=90;	data[28][9] <=61;	data[29][9] <=234;	data[30][9] <=25;	data[31][9] <=166;
    data[0][10] <=93;	data[1][10] <=114;	data[2][10] <=73;	data[3][10] <=130;	data[4][10] <=178;	data[5][10] <=11;	data[6][10] <=182;	data[7][10] <=149;	data[8][10] <=109;	data[9][10] <=50;	data[10][10] <=111;	data[11][10] <=230;	data[12][10] <=118;	data[13][10] <=135;	data[14][10] <=221;	data[15][10] <=161;	data[16][10] <=135;	data[17][10] <=219;	data[18][10] <=110;	data[19][10] <=136;	data[20][10] <=241;	data[21][10] <=250;	data[22][10] <=204;	data[23][10] <=41;	data[24][10] <=255;	data[25][10] <=118;	data[26][10] <=36;	data[27][10] <=116;	data[28][10] <=140;	data[29][10] <=216;	data[30][10] <=22;	data[31][10] <=173;
    data[0][11] <=23;	data[1][11] <=8;	data[2][11] <=239;	data[3][11] <=174;	data[4][11] <=140;	data[5][11] <=158;	data[6][11] <=134;	data[7][11] <=96;	data[8][11] <=141;	data[9][11] <=253;	data[10][11] <=212;	data[11][11] <=60;	data[12][11] <=253;	data[13][11] <=130;	data[14][11] <=65;	data[15][11] <=215;	data[16][11] <=108;	data[17][11] <=18;	data[18][11] <=160;	data[19][11] <=42;	data[20][11] <=43;	data[21][11] <=254;	data[22][11] <=22;	data[23][11] <=181;	data[24][11] <=123;	data[25][11] <=185;	data[26][11] <=222;	data[27][11] <=59;	data[28][11] <=231;	data[29][11] <=204;	data[30][11] <=151;	data[31][11] <=6;
    data[0][12] <=146;	data[1][12] <=195;	data[2][12] <=129;	data[3][12] <=135;	data[4][12] <=181;	data[5][12] <=29;	data[6][12] <=9;	data[7][12] <=161;	data[8][12] <=116;	data[9][12] <=47;	data[10][12] <=50;	data[11][12] <=189;	data[12][12] <=82;	data[13][12] <=157;	data[14][12] <=9;	data[15][12] <=71;	data[16][12] <=39;	data[17][12] <=192;	data[18][12] <=170;	data[19][12] <=145;	data[20][12] <=126;	data[21][12] <=151;	data[22][12] <=245;	data[23][12] <=30;	data[24][12] <=46;	data[25][12] <=236;	data[26][12] <=87;	data[27][12] <=78;	data[28][12] <=56;	data[29][12] <=25;	data[30][12] <=142;	data[31][12] <=129;
    data[0][13] <=234;	data[1][13] <=252;	data[2][13] <=5;	data[3][13] <=250;	data[4][13] <=211;	data[5][13] <=173;	data[6][13] <=175;	data[7][13] <=65;	data[8][13] <=247;	data[9][13] <=180;	data[10][13] <=178;	data[11][13] <=116;	data[12][13] <=155;	data[13][13] <=67;	data[14][13] <=36;	data[15][13] <=161;	data[16][13] <=158;	data[17][13] <=92;	data[18][13] <=177;	data[19][13] <=111;	data[20][13] <=57;	data[21][13] <=27;	data[22][13] <=183;	data[23][13] <=189;	data[24][13] <=125;	data[25][13] <=247;	data[26][13] <=40;	data[27][13] <=95;	data[28][13] <=84;	data[29][13] <=161;	data[30][13] <=41;	data[31][13] <=165;
    data[0][14] <=62;	data[1][14] <=177;	data[2][14] <=11;	data[3][14] <=237;	data[4][14] <=80;	data[5][14] <=79;	data[6][14] <=52;	data[7][14] <=44;	data[8][14] <=201;	data[9][14] <=159;	data[10][14] <=68;	data[11][14] <=240;	data[12][14] <=125;	data[13][14] <=222;	data[14][14] <=150;	data[15][14] <=160;	data[16][14] <=32;	data[17][14] <=246;	data[18][14] <=98;	data[19][14] <=59;	data[20][14] <=139;	data[21][14] <=27;	data[22][14] <=239;	data[23][14] <=249;	data[24][14] <=38;	data[25][14] <=140;	data[26][14] <=173;	data[27][14] <=35;	data[28][14] <=107;	data[29][14] <=200;	data[30][14] <=200;	data[31][14] <=21;
    data[0][15] <=225;	data[1][15] <=70;	data[2][15] <=239;	data[3][15] <=78;	data[4][15] <=241;	data[5][15] <=245;	data[6][15] <=19;	data[7][15] <=137;	data[8][15] <=10;	data[9][15] <=98;	data[10][15] <=91;	data[11][15] <=210;	data[12][15] <=17;	data[13][15] <=165;	data[14][15] <=6;	data[15][15] <=67;	data[16][15] <=227;	data[17][15] <=23;	data[18][15] <=3;	data[19][15] <=75;	data[20][15] <=167;	data[21][15] <=199;	data[22][15] <=120;	data[23][15] <=112;	data[24][15] <=59;	data[25][15] <=97;	data[26][15] <=143;	data[27][15] <=25;	data[28][15] <=22;	data[29][15] <=215;	data[30][15] <=67;	data[31][15] <=223;
	
	data[31][0] <=229;	data[32][0] <=82;	data[33][0] <=6;	data[34][0] <=247;	data[35][0] <=187;	data[36][0] <=155;	data[37][0] <=188;	data[38][0] <=132;	data[39][0] <=181;	data[40][0] <=129;	data[41][0] <=230;	data[42][0] <=236;	data[43][0] <=179;	data[44][0] <=172;	data[45][0] <=119;	data[46][0] <=194;	data[47][0] <=110;	data[48][0] <=201;	data[49][0] <=207;	data[50][0] <=16;	data[51][0] <=167;	data[52][0] <=187;	data[53][0] <=248;	data[54][0] <=152;	data[55][0] <=181;	data[56][0] <=71;	data[57][0] <=122;	data[58][0] <=178;	data[59][0] <=122;	data[60][0] <=57;	data[61][0] <=113;	data[62][0] <=106;	data[63][0] <=70;
    data[31][1] <=148;	data[32][1] <=30;	data[33][1] <=231;	data[34][1] <=211;	data[35][1] <=137;	data[36][1] <=28;	data[37][1] <=139;	data[38][1] <=128;	data[39][1] <=245;	data[40][1] <=193;	data[41][1] <=110;	data[42][1] <=135;	data[43][1] <=5;	data[44][1] <=198;	data[45][1] <=34;	data[46][1] <=193;	data[47][1] <=73;	data[48][1] <=44;	data[49][1] <=232;	data[50][1] <=167;	data[51][1] <=226;	data[52][1] <=30;	data[53][1] <=91;	data[54][1] <=163;	data[55][1] <=202;	data[56][1] <=86;	data[57][1] <=135;	data[58][1] <=123;	data[59][1] <=213;	data[60][1] <=241;	data[61][1] <=180;	data[62][1] <=192;	data[63][1] <=38;
    data[31][2] <=246;	data[32][2] <=193;	data[33][2] <=109;	data[34][2] <=69;	data[35][2] <=91;	data[36][2] <=244;	data[37][2] <=133;	data[38][2] <=132;	data[39][2] <=216;	data[40][2] <=231;	data[41][2] <=53;	data[42][2] <=226;	data[43][2] <=231;	data[44][2] <=3;	data[45][2] <=54;	data[46][2] <=15;	data[47][2] <=135;	data[48][2] <=110;	data[49][2] <=57;	data[50][2] <=20;	data[51][2] <=40;	data[52][2] <=201;	data[53][2] <=238;	data[54][2] <=16;	data[55][2] <=156;	data[56][2] <=2;	data[57][2] <=80;	data[58][2] <=28;	data[59][2] <=238;	data[60][2] <=99;	data[61][2] <=168;	data[62][2] <=23;	data[63][2] <=126;
    data[31][3] <=56;	data[32][3] <=127;	data[33][3] <=195;	data[34][3] <=151;	data[35][3] <=138;	data[36][3] <=150;	data[37][3] <=84;	data[38][3] <=143;	data[39][3] <=133;	data[40][3] <=65;	data[41][3] <=84;	data[42][3] <=221;	data[43][3] <=55;	data[44][3] <=78;	data[45][3] <=9;	data[46][3] <=138;	data[47][3] <=25;	data[48][3] <=176;	data[49][3] <=2;	data[50][3] <=91;	data[51][3] <=251;	data[52][3] <=18;	data[53][3] <=197;	data[54][3] <=83;	data[55][3] <=168;	data[56][3] <=4;	data[57][3] <=191;	data[58][3] <=104;	data[59][3] <=151;	data[60][3] <=201;	data[61][3] <=225;	data[62][3] <=207;	data[63][3] <=219;
    data[31][4] <=159;	data[32][4] <=195;	data[33][4] <=146;	data[34][4] <=85;	data[35][4] <=18;	data[36][4] <=127;	data[37][4] <=172;	data[38][4] <=234;	data[39][4] <=12;	data[40][4] <=107;	data[41][4] <=4;	data[42][4] <=186;	data[43][4] <=100;	data[44][4] <=238;	data[45][4] <=188;	data[46][4] <=222;	data[47][4] <=231;	data[48][4] <=15;	data[49][4] <=95;	data[50][4] <=222;	data[51][4] <=20;	data[52][4] <=2;	data[53][4] <=10;	data[54][4] <=176;	data[55][4] <=103;	data[56][4] <=46;	data[57][4] <=72;	data[58][4] <=222;	data[59][4] <=114;	data[60][4] <=240;	data[61][4] <=229;	data[62][4] <=169;	data[63][4] <=24;
    data[31][5] <=233;	data[32][5] <=253;	data[33][5] <=15;	data[34][5] <=15;	data[35][5] <=230;	data[36][5] <=117;	data[37][5] <=10;	data[38][5] <=248;	data[39][5] <=186;	data[40][5] <=218;	data[41][5] <=63;	data[42][5] <=87;	data[43][5] <=124;	data[44][5] <=248;	data[45][5] <=27;	data[46][5] <=127;	data[47][5] <=76;	data[48][5] <=108;	data[49][5] <=205;	data[50][5] <=241;	data[51][5] <=80;	data[52][5] <=220;	data[53][5] <=218;	data[54][5] <=253;	data[55][5] <=14;	data[56][5] <=215;	data[57][5] <=17;	data[58][5] <=110;	data[59][5] <=222;	data[60][5] <=46;	data[61][5] <=208;	data[62][5] <=36;	data[63][5] <=240;
    data[31][6] <=156;	data[32][6] <=48;	data[33][6] <=160;	data[34][6] <=130;	data[35][6] <=95;	data[36][6] <=173;	data[37][6] <=246;	data[38][6] <=210;	data[39][6] <=75;	data[40][6] <=183;	data[41][6] <=114;	data[42][6] <=186;	data[43][6] <=161;	data[44][6] <=146;	data[45][6] <=127;	data[46][6] <=218;	data[47][6] <=150;	data[48][6] <=169;	data[49][6] <=104;	data[50][6] <=117;	data[51][6] <=120;	data[52][6] <=41;	data[53][6] <=154;	data[54][6] <=127;	data[55][6] <=131;	data[56][6] <=152;	data[57][6] <=57;	data[58][6] <=213;	data[59][6] <=176;	data[60][6] <=44;	data[61][6] <=180;	data[62][6] <=156;	data[63][6] <=18;
    data[31][7] <=192;	data[32][7] <=245;	data[33][7] <=77;	data[34][7] <=64;	data[35][7] <=64;	data[36][7] <=29;	data[37][7] <=30;	data[38][7] <=15;	data[39][7] <=67;	data[40][7] <=113;	data[41][7] <=62;	data[42][7] <=62;	data[43][7] <=115;	data[44][7] <=163;	data[45][7] <=38;	data[46][7] <=181;	data[47][7] <=235;	data[48][7] <=201;	data[49][7] <=250;	data[50][7] <=45;	data[51][7] <=250;	data[52][7] <=139;	data[53][7] <=185;	data[54][7] <=33;	data[55][7] <=90;	data[56][7] <=70;	data[57][7] <=7;	data[58][7] <=92;	data[59][7] <=137;	data[60][7] <=240;	data[61][7] <=210;	data[62][7] <=52;	data[63][7] <=166;
    data[31][8] <=33;	data[32][8] <=252;	data[33][8] <=55;	data[34][8] <=125;	data[35][8] <=214;	data[36][8] <=2;	data[37][8] <=85;	data[38][8] <=63;	data[39][8] <=169;	data[40][8] <=17;	data[41][8] <=62;	data[42][8] <=157;	data[43][8] <=122;	data[44][8] <=18;	data[45][8] <=255;	data[46][8] <=138;	data[47][8] <=52;	data[48][8] <=210;	data[49][8] <=254;	data[50][8] <=68;	data[51][8] <=182;	data[52][8] <=24;	data[53][8] <=178;	data[54][8] <=208;	data[55][8] <=12;	data[56][8] <=217;	data[57][8] <=237;	data[58][8] <=128;	data[59][8] <=60;	data[60][8] <=172;	data[61][8] <=83;	data[62][8] <=247;	data[63][8] <=237;
    data[31][9] <=166;	data[32][9] <=186;	data[33][9] <=138;	data[34][9] <=237;	data[35][9] <=78;	data[36][9] <=224;	data[37][9] <=251;	data[38][9] <=235;	data[39][9] <=133;	data[40][9] <=96;	data[41][9] <=156;	data[42][9] <=56;	data[43][9] <=176;	data[44][9] <=125;	data[45][9] <=99;	data[46][9] <=43;	data[47][9] <=142;	data[48][9] <=165;	data[49][9] <=33;	data[50][9] <=249;	data[51][9] <=88;	data[52][9] <=163;	data[53][9] <=158;	data[54][9] <=1;	data[55][9] <=152;	data[56][9] <=122;	data[57][9] <=209;	data[58][9] <=112;	data[59][9] <=163;	data[60][9] <=224;	data[61][9] <=246;	data[62][9] <=97;	data[63][9] <=3;
    data[31][10] <=173;	data[32][10] <=104;	data[33][10] <=119;	data[34][10] <=129;	data[35][10] <=1;	data[36][10] <=104;	data[37][10] <=86;	data[38][10] <=212;	data[39][10] <=246;	data[40][10] <=233;	data[41][10] <=164;	data[42][10] <=255;	data[43][10] <=41;	data[44][10] <=200;	data[45][10] <=23;	data[46][10] <=136;	data[47][10] <=213;	data[48][10] <=213;	data[49][10] <=46;	data[50][10] <=231;	data[51][10] <=70;	data[52][10] <=109;	data[53][10] <=84;	data[54][10] <=219;	data[55][10] <=8;	data[56][10] <=185;	data[57][10] <=14;	data[58][10] <=207;	data[59][10] <=86;	data[60][10] <=76;	data[61][10] <=18;	data[62][10] <=116;	data[63][10] <=221;
    data[31][11] <=6;	data[32][11] <=166;	data[33][11] <=108;	data[34][11] <=21;	data[35][11] <=130;	data[36][11] <=239;	data[37][11] <=177;	data[38][11] <=252;	data[39][11] <=111;	data[40][11] <=73;	data[41][11] <=248;	data[42][11] <=62;	data[43][11] <=9;	data[44][11] <=215;	data[45][11] <=174;	data[46][11] <=53;	data[47][11] <=28;	data[48][11] <=62;	data[49][11] <=65;	data[50][11] <=150;	data[51][11] <=153;	data[52][11] <=72;	data[53][11] <=226;	data[54][11] <=183;	data[55][11] <=33;	data[56][11] <=217;	data[57][11] <=16;	data[58][11] <=15;	data[59][11] <=214;	data[60][11] <=232;	data[61][11] <=39;	data[62][11] <=5;	data[63][11] <=118;
    data[31][12] <=129;	data[32][12] <=160;	data[33][12] <=111;	data[34][12] <=79;	data[35][12] <=31;	data[36][12] <=204;	data[37][12] <=180;	data[38][12] <=24;	data[39][12] <=245;	data[40][12] <=236;	data[41][12] <=36;	data[42][12] <=254;	data[43][12] <=34;	data[44][12] <=35;	data[45][12] <=150;	data[46][12] <=237;	data[47][12] <=255;	data[48][12] <=154;	data[49][12] <=202;	data[50][12] <=226;	data[51][12] <=228;	data[52][12] <=171;	data[53][12] <=104;	data[54][12] <=235;	data[55][12] <=168;	data[56][12] <=23;	data[57][12] <=161;	data[58][12] <=137;	data[59][12] <=133;	data[60][12] <=19;	data[61][12] <=194;	data[62][12] <=232;	data[63][12] <=152;
    data[31][13] <=165;	data[32][13] <=234;	data[33][13] <=223;	data[34][13] <=235;	data[35][13] <=121;	data[36][13] <=122;	data[37][13] <=177;	data[38][13] <=132;	data[39][13] <=0;	data[40][13] <=231;	data[41][13] <=23;	data[42][13] <=172;	data[43][13] <=186;	data[44][13] <=225;	data[45][13] <=87;	data[46][13] <=18;	data[47][13] <=255;	data[48][13] <=15;	data[49][13] <=177;	data[50][13] <=22;	data[51][13] <=59;	data[52][13] <=85;	data[53][13] <=208;	data[54][13] <=241;	data[55][13] <=244;	data[56][13] <=33;	data[57][13] <=10;	data[58][13] <=12;	data[59][13] <=222;	data[60][13] <=165;	data[61][13] <=157;	data[62][13] <=173;	data[63][13] <=72;
    data[31][14] <=21;	data[32][14] <=3;	data[33][14] <=29;	data[34][14] <=148;	data[35][14] <=151;	data[36][14] <=231;	data[37][14] <=33;	data[38][14] <=51;	data[39][14] <=181;	data[40][14] <=59;	data[41][14] <=49;	data[42][14] <=223;	data[43][14] <=27;	data[44][14] <=147;	data[45][14] <=210;	data[46][14] <=66;	data[47][14] <=108;	data[48][14] <=36;	data[49][14] <=212;	data[50][14] <=24;	data[51][14] <=219;	data[52][14] <=3;	data[53][14] <=17;	data[54][14] <=234;	data[55][14] <=144;	data[56][14] <=146;	data[57][14] <=219;	data[58][14] <=20;	data[59][14] <=42;	data[60][14] <=116;	data[61][14] <=158;	data[62][14] <=127;	data[63][14] <=13;
    data[31][15] <=223;	data[32][15] <=250;	data[33][15] <=131;	data[34][15] <=125;	data[35][15] <=162;	data[36][15] <=207;	data[37][15] <=196;	data[38][15] <=29;	data[39][15] <=150;	data[40][15] <=233;	data[41][15] <=114;	data[42][15] <=67;	data[43][15] <=116;	data[44][15] <=36;	data[45][15] <=184;	data[46][15] <=3;	data[47][15] <=197;	data[48][15] <=67;	data[49][15] <=209;	data[50][15] <=21;	data[51][15] <=72;	data[52][15] <=4;	data[53][15] <=59;	data[54][15] <=169;	data[55][15] <=232;	data[56][15] <=200;	data[57][15] <=80;	data[58][15] <=158;	data[59][15] <=239;	data[60][15] <=236;	data[61][15] <=104;	data[62][15] <=60;	data[63][15] <=33;

	data[64][0] <=249;	data[65][0] <=48;	data[66][0] <=84;	data[67][0] <=91;	data[68][0] <=125;	data[69][0] <=85;	data[70][0] <=98;	data[71][0] <=215;	data[72][0] <=166;	data[73][0] <=11;	data[74][0] <=33;	data[75][0] <=241;	data[76][0] <=210;	data[77][0] <=49;	data[78][0] <=15;	data[79][0] <=184;	data[80][0] <=66;	data[81][0] <=160;	data[82][0] <=30;	data[83][0] <=59;	data[84][0] <=68;	data[85][0] <=142;	data[86][0] <=34;	data[87][0] <=67;	data[88][0] <=248;	data[89][0] <=66;	data[90][0] <=106;	data[91][0] <=79;	data[92][0] <=235;	data[93][0] <=169;	data[94][0] <=218;	data[95][0] <=138;	data[96][0] <=129;	data[97][0] <=220;	data[98][0] <=49;	data[99][0] <=239;	data[100][0] <=146;	data[101][0] <=75;	data[102][0] <=196;	data[103][0] <=132;	data[104][0] <=206;	data[105][0] <=85;	data[106][0] <=182;	data[107][0] <=178;	data[108][0] <=175;	data[109][0] <=34;	data[110][0] <=234;	data[111][0] <=194;	data[112][0] <=63;	data[113][0] <=108;	data[114][0] <=87;	data[115][0] <=65;	data[116][0] <=212;	data[117][0] <=195;	data[118][0] <=128;	data[119][0] <=188;	data[120][0] <=27;	data[121][0] <=155;	data[122][0] <=12;	data[123][0] <=53;	data[124][0] <=126;	data[125][0] <=67;	data[126][0] <=231;	data[127][0] <=124;
	data[64][1] <=98;	data[65][1] <=14;	data[66][1] <=246;	data[67][1] <=193;	data[68][1] <=96;	data[69][1] <=113;	data[70][1] <=115;	data[71][1] <=121;	data[72][1] <=217;	data[73][1] <=247;	data[74][1] <=220;	data[75][1] <=50;	data[76][1] <=81;	data[77][1] <=134;	data[78][1] <=57;	data[79][1] <=63;	data[80][1] <=177;	data[81][1] <=116;	data[82][1] <=152;	data[83][1] <=225;	data[84][1] <=113;	data[85][1] <=178;	data[86][1] <=240;	data[87][1] <=48;	data[88][1] <=199;	data[89][1] <=6;	data[90][1] <=28;	data[91][1] <=29;	data[92][1] <=172;	data[93][1] <=186;	data[94][1] <=227;	data[95][1] <=44;	data[96][1] <=27;	data[97][1] <=67;	data[98][1] <=25;	data[99][1] <=90;	data[100][1] <=249;	data[101][1] <=106;	data[102][1] <=6;	data[103][1] <=145;	data[104][1] <=26;	data[105][1] <=178;	data[106][1] <=61;	data[107][1] <=88;	data[108][1] <=141;	data[109][1] <=237;	data[110][1] <=34;	data[111][1] <=251;	data[112][1] <=21;	data[113][1] <=199;	data[114][1] <=244;	data[115][1] <=18;	data[116][1] <=162;	data[117][1] <=56;	data[118][1] <=21;	data[119][1] <=4;	data[120][1] <=156;	data[121][1] <=67;	data[122][1] <=3;	data[123][1] <=249;	data[124][1] <=174;	data[125][1] <=12;	data[126][1] <=96;	data[127][1] <=81;
	data[64][2] <=236;	data[65][2] <=65;	data[66][2] <=184;	data[67][2] <=11;	data[68][2] <=149;	data[69][2] <=89;	data[70][2] <=25;	data[71][2] <=152;	data[72][2] <=123;	data[73][2] <=246;	data[74][2] <=101;	data[75][2] <=113;	data[76][2] <=57;	data[77][2] <=55;	data[78][2] <=129;	data[79][2] <=43;	data[80][2] <=69;	data[81][2] <=79;	data[82][2] <=15;	data[83][2] <=48;	data[84][2] <=17;	data[85][2] <=236;	data[86][2] <=173;	data[87][2] <=184;	data[88][2] <=194;	data[89][2] <=110;	data[90][2] <=8;	data[91][2] <=112;	data[92][2] <=63;	data[93][2] <=82;	data[94][2] <=33;	data[95][2] <=71;	data[96][2] <=239;	data[97][2] <=218;	data[98][2] <=36;	data[99][2] <=93;	data[100][2] <=170;	data[101][2] <=199;	data[102][2] <=157;	data[103][2] <=236;	data[104][2] <=130;	data[105][2] <=20;	data[106][2] <=19;	data[107][2] <=45;	data[108][2] <=211;	data[109][2] <=43;	data[110][2] <=252;	data[111][2] <=234;	data[112][2] <=185;	data[113][2] <=199;	data[114][2] <=51;	data[115][2] <=45;	data[116][2] <=107;	data[117][2] <=202;	data[118][2] <=243;	data[119][2] <=216;	data[120][2] <=154;	data[121][2] <=75;	data[122][2] <=52;	data[123][2] <=30;	data[124][2] <=130;	data[125][2] <=253;	data[126][2] <=174;	data[127][2] <=170;
	data[64][3] <=247;	data[65][3] <=174;	data[66][3] <=6;	data[67][3] <=8;	data[68][3] <=148;	data[69][3] <=31;	data[70][3] <=125;	data[71][3] <=204;	data[72][3] <=29;	data[73][3] <=23;	data[74][3] <=221;	data[75][3] <=185;	data[76][3] <=254;	data[77][3] <=104;	data[78][3] <=30;	data[79][3] <=93;	data[80][3] <=200;	data[81][3] <=102;	data[82][3] <=192;	data[83][3] <=99;	data[84][3] <=176;	data[85][3] <=15;	data[86][3] <=187;	data[87][3] <=247;	data[88][3] <=206;	data[89][3] <=91;	data[90][3] <=255;	data[91][3] <=106;	data[92][3] <=164;	data[93][3] <=179;	data[94][3] <=189;	data[95][3] <=134;	data[96][3] <=241;	data[97][3] <=165;	data[98][3] <=169;	data[99][3] <=56;	data[100][3] <=157;	data[101][3] <=120;	data[102][3] <=101;	data[103][3] <=55;	data[104][3] <=70;	data[105][3] <=130;	data[106][3] <=189;	data[107][3] <=59;	data[108][3] <=211;	data[109][3] <=95;	data[110][3] <=158;	data[111][3] <=217;	data[112][3] <=13;	data[113][3] <=7;	data[114][3] <=207;	data[115][3] <=221;	data[116][3] <=51;	data[117][3] <=52;	data[118][3] <=191;	data[119][3] <=38;	data[120][3] <=197;	data[121][3] <=83;	data[122][3] <=154;	data[123][3] <=69;	data[124][3] <=29;	data[125][3] <=68;	data[126][3] <=131;	data[127][3] <=28;
	data[64][4] <=147;	data[65][4] <=173;	data[66][4] <=26;	data[67][4] <=237;	data[68][4] <=45;	data[69][4] <=35;	data[70][4] <=141;	data[71][4] <=126;	data[72][4] <=178;	data[73][4] <=69;	data[74][4] <=252;	data[75][4] <=115;	data[76][4] <=15;	data[77][4] <=121;	data[78][4] <=64;	data[79][4] <=32;	data[80][4] <=89;	data[81][4] <=147;	data[82][4] <=189;	data[83][4] <=166;	data[84][4] <=139;	data[85][4] <=209;	data[86][4] <=121;	data[87][4] <=90;	data[88][4] <=173;	data[89][4] <=56;	data[90][4] <=139;	data[91][4] <=247;	data[92][4] <=12;	data[93][4] <=72;	data[94][4] <=211;	data[95][4] <=82;	data[96][4] <=254;	data[97][4] <=185;	data[98][4] <=186;	data[99][4] <=196;	data[100][4] <=171;	data[101][4] <=240;	data[102][4] <=186;	data[103][4] <=128;	data[104][4] <=111;	data[105][4] <=142;	data[106][4] <=6;	data[107][4] <=21;	data[108][4] <=73;	data[109][4] <=110;	data[110][4] <=217;	data[111][4] <=78;	data[112][4] <=88;	data[113][4] <=98;	data[114][4] <=153;	data[115][4] <=162;	data[116][4] <=245;	data[117][4] <=194;	data[118][4] <=16;	data[119][4] <=136;	data[120][4] <=203;	data[121][4] <=237;	data[122][4] <=0;	data[123][4] <=16;	data[124][4] <=81;	data[125][4] <=26;	data[126][4] <=115;	data[127][4] <=100;
	data[64][5] <=119;	data[65][5] <=154;	data[66][5] <=155;	data[67][5] <=79;	data[68][5] <=161;	data[69][5] <=151;	data[70][5] <=120;	data[71][5] <=25;	data[72][5] <=97;	data[73][5] <=237;	data[74][5] <=76;	data[75][5] <=104;	data[76][5] <=101;	data[77][5] <=27;	data[78][5] <=165;	data[79][5] <=44;	data[80][5] <=102;	data[81][5] <=126;	data[82][5] <=116;	data[83][5] <=87;	data[84][5] <=240;	data[85][5] <=34;	data[86][5] <=24;	data[87][5] <=246;	data[88][5] <=208;	data[89][5] <=58;	data[90][5] <=177;	data[91][5] <=80;	data[92][5] <=30;	data[93][5] <=180;	data[94][5] <=110;	data[95][5] <=3;	data[96][5] <=20;	data[97][5] <=133;	data[98][5] <=155;	data[99][5] <=41;	data[100][5] <=58;	data[101][5] <=249;	data[102][5] <=139;	data[103][5] <=56;	data[104][5] <=91;	data[105][5] <=201;	data[106][5] <=40;	data[107][5] <=4;	data[108][5] <=50;	data[109][5] <=211;	data[110][5] <=243;	data[111][5] <=227;	data[112][5] <=111;	data[113][5] <=21;	data[114][5] <=39;	data[115][5] <=199;	data[116][5] <=161;	data[117][5] <=121;	data[118][5] <=113;	data[119][5] <=117;	data[120][5] <=242;	data[121][5] <=225;	data[122][5] <=190;	data[123][5] <=228;	data[124][5] <=37;	data[125][5] <=217;	data[126][5] <=86;	data[127][5] <=95;
	data[64][6] <=139;	data[65][6] <=196;	data[66][6] <=227;	data[67][6] <=56;	data[68][6] <=253;	data[69][6] <=236;	data[70][6] <=208;	data[71][6] <=146;	data[72][6] <=76;	data[73][6] <=116;	data[74][6] <=14;	data[75][6] <=70;	data[76][6] <=76;	data[77][6] <=15;	data[78][6] <=94;	data[79][6] <=75;	data[80][6] <=167;	data[81][6] <=159;	data[82][6] <=51;	data[83][6] <=75;	data[84][6] <=118;	data[85][6] <=115;	data[86][6] <=209;	data[87][6] <=175;	data[88][6] <=169;	data[89][6] <=233;	data[90][6] <=20;	data[91][6] <=220;	data[92][6] <=143;	data[93][6] <=162;	data[94][6] <=75;	data[95][6] <=21;	data[96][6] <=201;	data[97][6] <=184;	data[98][6] <=200;	data[99][6] <=180;	data[100][6] <=195;	data[101][6] <=205;	data[102][6] <=86;	data[103][6] <=82;	data[104][6] <=218;	data[105][6] <=133;	data[106][6] <=81;	data[107][6] <=92;	data[108][6] <=124;	data[109][6] <=56;	data[110][6] <=82;	data[111][6] <=5;	data[112][6] <=43;	data[113][6] <=5;	data[114][6] <=132;	data[115][6] <=30;	data[116][6] <=230;	data[117][6] <=122;	data[118][6] <=40;	data[119][6] <=244;	data[120][6] <=39;	data[121][6] <=182;	data[122][6] <=246;	data[123][6] <=208;	data[124][6] <=221;	data[125][6] <=129;	data[126][6] <=217;	data[127][6] <=66;
	data[64][7] <=172;	data[65][7] <=200;	data[66][7] <=214;	data[67][7] <=176;	data[68][7] <=191;	data[69][7] <=188;	data[70][7] <=84;	data[71][7] <=144;	data[72][7] <=147;	data[73][7] <=11;	data[74][7] <=186;	data[75][7] <=84;	data[76][7] <=31;	data[77][7] <=59;	data[78][7] <=143;	data[79][7] <=114;	data[80][7] <=104;	data[81][7] <=117;	data[82][7] <=252;	data[83][7] <=230;	data[84][7] <=88;	data[85][7] <=241;	data[86][7] <=35;	data[87][7] <=186;	data[88][7] <=118;	data[89][7] <=58;	data[90][7] <=192;	data[91][7] <=1;	data[92][7] <=96;	data[93][7] <=203;	data[94][7] <=161;	data[95][7] <=172;	data[96][7] <=140;	data[97][7] <=154;	data[98][7] <=129;	data[99][7] <=53;	data[100][7] <=98;	data[101][7] <=94;	data[102][7] <=91;	data[103][7] <=37;	data[104][7] <=106;	data[105][7] <=169;	data[106][7] <=58;	data[107][7] <=63;	data[108][7] <=109;	data[109][7] <=16;	data[110][7] <=51;	data[111][7] <=226;	data[112][7] <=146;	data[113][7] <=235;	data[114][7] <=106;	data[115][7] <=121;	data[116][7] <=19;	data[117][7] <=87;	data[118][7] <=200;	data[119][7] <=84;	data[120][7] <=250;	data[121][7] <=200;	data[122][7] <=64;	data[123][7] <=230;	data[124][7] <=219;	data[125][7] <=241;	data[126][7] <=255;	data[127][7] <=195;
	data[64][8] <=9;	data[65][8] <=42;	data[66][8] <=88;	data[67][8] <=35;	data[68][8] <=66;	data[69][8] <=141;	data[70][8] <=233;	data[71][8] <=34;	data[72][8] <=7;	data[73][8] <=249;	data[74][8] <=33;	data[75][8] <=204;	data[76][8] <=73;	data[77][8] <=131;	data[78][8] <=189;	data[79][8] <=125;	data[80][8] <=7;	data[81][8] <=60;	data[82][8] <=133;	data[83][8] <=113;	data[84][8] <=7;	data[85][8] <=230;	data[86][8] <=160;	data[87][8] <=227;	data[88][8] <=240;	data[89][8] <=62;	data[90][8] <=223;	data[91][8] <=13;	data[92][8] <=72;	data[93][8] <=164;	data[94][8] <=88;	data[95][8] <=43;	data[96][8] <=251;	data[97][8] <=67;	data[98][8] <=24;	data[99][8] <=184;	data[100][8] <=165;	data[101][8] <=146;	data[102][8] <=247;	data[103][8] <=90;	data[104][8] <=54;	data[105][8] <=2;	data[106][8] <=165;	data[107][8] <=210;	data[108][8] <=82;	data[109][8] <=128;	data[110][8] <=255;	data[111][8] <=234;	data[112][8] <=176;	data[113][8] <=100;	data[114][8] <=182;	data[115][8] <=63;	data[116][8] <=219;	data[117][8] <=23;	data[118][8] <=51;	data[119][8] <=54;	data[120][8] <=103;	data[121][8] <=7;	data[122][8] <=38;	data[123][8] <=37;	data[124][8] <=222;	data[125][8] <=166;	data[126][8] <=48;	data[127][8] <=33;
	data[64][9] <=49;	data[65][9] <=76;	data[66][9] <=125;	data[67][9] <=239;	data[68][9] <=136;	data[69][9] <=192;	data[70][9] <=82;	data[71][9] <=141;	data[72][9] <=210;	data[73][9] <=252;	data[74][9] <=203;	data[75][9] <=153;	data[76][9] <=173;	data[77][9] <=190;	data[78][9] <=182;	data[79][9] <=160;	data[80][9] <=57;	data[81][9] <=133;	data[82][9] <=220;	data[83][9] <=191;	data[84][9] <=56;	data[85][9] <=38;	data[86][9] <=180;	data[87][9] <=209;	data[88][9] <=108;	data[89][9] <=197;	data[90][9] <=76;	data[91][9] <=106;	data[92][9] <=201;	data[93][9] <=80;	data[94][9] <=230;	data[95][9] <=192;	data[96][9] <=99;	data[97][9] <=235;	data[98][9] <=223;	data[99][9] <=162;	data[100][9] <=98;	data[101][9] <=95;	data[102][9] <=93;	data[103][9] <=109;	data[104][9] <=23;	data[105][9] <=78;	data[106][9] <=196;	data[107][9] <=213;	data[108][9] <=109;	data[109][9] <=93;	data[110][9] <=250;	data[111][9] <=142;	data[112][9] <=69;	data[113][9] <=111;	data[114][9] <=172;	data[115][9] <=68;	data[116][9] <=246;	data[117][9] <=197;	data[118][9] <=5;	data[119][9] <=20;	data[120][9] <=104;	data[121][9] <=198;	data[122][9] <=239;	data[123][9] <=169;	data[124][9] <=96;	data[125][9] <=87;	data[126][9] <=29;	data[127][9] <=164;
	data[64][10] <=146;	data[65][10] <=115;	data[66][10] <=62;	data[67][10] <=105;	data[68][10] <=92;	data[69][10] <=96;	data[70][10] <=11;	data[71][10] <=72;	data[72][10] <=61;	data[73][10] <=127;	data[74][10] <=94;	data[75][10] <=145;	data[76][10] <=42;	data[77][10] <=107;	data[78][10] <=56;	data[79][10] <=16;	data[80][10] <=84;	data[81][10] <=169;	data[82][10] <=46;	data[83][10] <=86;	data[84][10] <=226;	data[85][10] <=152;	data[86][10] <=29;	data[87][10] <=229;	data[88][10] <=246;	data[89][10] <=29;	data[90][10] <=152;	data[91][10] <=175;	data[92][10] <=212;	data[93][10] <=184;	data[94][10] <=253;	data[95][10] <=232;	data[96][10] <=64;	data[97][10] <=102;	data[98][10] <=164;	data[99][10] <=158;	data[100][10] <=244;	data[101][10] <=159;	data[102][10] <=105;	data[103][10] <=27;	data[104][10] <=66;	data[105][10] <=125;	data[106][10] <=41;	data[107][10] <=225;	data[108][10] <=180;	data[109][10] <=190;	data[110][10] <=253;	data[111][10] <=88;	data[112][10] <=218;	data[113][10] <=204;	data[114][10] <=164;	data[115][10] <=251;	data[116][10] <=135;	data[117][10] <=15;	data[118][10] <=150;	data[119][10] <=10;	data[120][10] <=50;	data[121][10] <=165;	data[122][10] <=82;	data[123][10] <=9;	data[124][10] <=196;	data[125][10] <=101;	data[126][10] <=94;	data[127][10] <=243;
	data[64][11] <=47;	data[65][11] <=186;	data[66][11] <=251;	data[67][11] <=28;	data[68][11] <=66;	data[69][11] <=62;	data[70][11] <=67;	data[71][11] <=33;	data[72][11] <=187;	data[73][11] <=4;	data[74][11] <=51;	data[75][11] <=210;	data[76][11] <=222;	data[77][11] <=183;	data[78][11] <=223;	data[79][11] <=87;	data[80][11] <=210;	data[81][11] <=51;	data[82][11] <=93;	data[83][11] <=51;	data[84][11] <=116;	data[85][11] <=7;	data[86][11] <=206;	data[87][11] <=128;	data[88][11] <=161;	data[89][11] <=242;	data[90][11] <=23;	data[91][11] <=219;	data[92][11] <=16;	data[93][11] <=42;	data[94][11] <=71;	data[95][11] <=133;	data[96][11] <=166;	data[97][11] <=109;	data[98][11] <=111;	data[99][11] <=25;	data[100][11] <=242;	data[101][11] <=92;	data[102][11] <=131;	data[103][11] <=230;	data[104][11] <=206;	data[105][11] <=199;	data[106][11] <=142;	data[107][11] <=73;	data[108][11] <=174;	data[109][11] <=73;	data[110][11] <=140;	data[111][11] <=159;	data[112][11] <=117;	data[113][11] <=202;	data[114][11] <=130;	data[115][11] <=216;	data[116][11] <=28;	data[117][11] <=108;	data[118][11] <=86;	data[119][11] <=164;	data[120][11] <=152;	data[121][11] <=52;	data[122][11] <=182;	data[123][11] <=138;	data[124][11] <=191;	data[125][11] <=203;	data[126][11] <=206;	data[127][11] <=53;
	data[64][12] <=62;	data[65][12] <=234;	data[66][12] <=17;	data[67][12] <=222;	data[68][12] <=32;	data[69][12] <=114;	data[70][12] <=188;	data[71][12] <=147;	data[72][12] <=193;	data[73][12] <=198;	data[74][12] <=30;	data[75][12] <=225;	data[76][12] <=51;	data[77][12] <=45;	data[78][12] <=160;	data[79][12] <=73;	data[80][12] <=143;	data[81][12] <=151;	data[82][12] <=75;	data[83][12] <=12;	data[84][12] <=53;	data[85][12] <=1;	data[86][12] <=46;	data[87][12] <=153;	data[88][12] <=8;	data[89][12] <=141;	data[90][12] <=10;	data[91][12] <=24;	data[92][12] <=105;	data[93][12] <=211;	data[94][12] <=149;	data[95][12] <=141;	data[96][12] <=35;	data[97][12] <=137;	data[98][12] <=95;	data[99][12] <=247;	data[100][12] <=120;	data[101][12] <=69;	data[102][12] <=46;	data[103][12] <=182;	data[104][12] <=126;	data[105][12] <=170;	data[106][12] <=241;	data[107][12] <=12;	data[108][12] <=58;	data[109][12] <=204;	data[110][12] <=243;	data[111][12] <=172;	data[112][12] <=207;	data[113][12] <=246;	data[114][12] <=6;	data[115][12] <=225;	data[116][12] <=124;	data[117][12] <=38;	data[118][12] <=159;	data[119][12] <=159;	data[120][12] <=73;	data[121][12] <=131;	data[122][12] <=77;	data[123][12] <=63;	data[124][12] <=250;	data[125][12] <=218;	data[126][12] <=101;	data[127][12] <=14;
	data[64][13] <=183;	data[65][13] <=212;	data[66][13] <=106;	data[67][13] <=178;	data[68][13] <=156;	data[69][13] <=243;	data[70][13] <=73;	data[71][13] <=173;	data[72][13] <=58;	data[73][13] <=50;	data[74][13] <=17;	data[75][13] <=104;	data[76][13] <=236;	data[77][13] <=192;	data[78][13] <=75;	data[79][13] <=160;	data[80][13] <=221;	data[81][13] <=225;	data[82][13] <=88;	data[83][13] <=243;	data[84][13] <=111;	data[85][13] <=162;	data[86][13] <=151;	data[87][13] <=239;	data[88][13] <=90;	data[89][13] <=93;	data[90][13] <=220;	data[91][13] <=136;	data[92][13] <=95;	data[93][13] <=241;	data[94][13] <=91;	data[95][13] <=115;	data[96][13] <=15;	data[97][13] <=172;	data[98][13] <=220;	data[99][13] <=122;	data[100][13] <=144;	data[101][13] <=75;	data[102][13] <=165;	data[103][13] <=121;	data[104][13] <=97;	data[105][13] <=251;	data[106][13] <=174;	data[107][13] <=127;	data[108][13] <=184;	data[109][13] <=254;	data[110][13] <=19;	data[111][13] <=192;	data[112][13] <=65;	data[113][13] <=92;	data[114][13] <=123;	data[115][13] <=80;	data[116][13] <=219;	data[117][13] <=188;	data[118][13] <=231;	data[119][13] <=165;	data[120][13] <=210;	data[121][13] <=152;	data[122][13] <=118;	data[123][13] <=2;	data[124][13] <=117;	data[125][13] <=160;	data[126][13] <=160;	data[127][13] <=159;
	data[64][14] <=27;	data[65][14] <=187;	data[66][14] <=136;	data[67][14] <=92;	data[68][14] <=89;	data[69][14] <=9;	data[70][14] <=146;	data[71][14] <=29;	data[72][14] <=164;	data[73][14] <=26;	data[74][14] <=123;	data[75][14] <=53;	data[76][14] <=128;	data[77][14] <=80;	data[78][14] <=51;	data[79][14] <=210;	data[80][14] <=64;	data[81][14] <=225;	data[82][14] <=99;	data[83][14] <=116;	data[84][14] <=20;	data[85][14] <=40;	data[86][14] <=231;	data[87][14] <=13;	data[88][14] <=132;	data[89][14] <=196;	data[90][14] <=12;	data[91][14] <=63;	data[92][14] <=140;	data[93][14] <=103;	data[94][14] <=195;	data[95][14] <=88;	data[96][14] <=255;	data[97][14] <=249;	data[98][14] <=17;	data[99][14] <=32;	data[100][14] <=228;	data[101][14] <=46;	data[102][14] <=163;	data[103][14] <=66;	data[104][14] <=255;	data[105][14] <=91;	data[106][14] <=236;	data[107][14] <=83;	data[108][14] <=4;	data[109][14] <=183;	data[110][14] <=121;	data[111][14] <=88;	data[112][14] <=49;	data[113][14] <=126;	data[114][14] <=210;	data[115][14] <=202;	data[116][14] <=41;	data[117][14] <=252;	data[118][14] <=179;	data[119][14] <=139;	data[120][14] <=169;	data[121][14] <=121;	data[122][14] <=117;	data[123][14] <=19;	data[124][14] <=254;	data[125][14] <=81;	data[126][14] <=94;	data[127][14] <=101;
	data[64][15] <=127;	data[65][15] <=172;	data[66][15] <=125;	data[67][15] <=23;	data[68][15] <=171;	data[69][15] <=200;	data[70][15] <=46;	data[71][15] <=201;	data[72][15] <=161;	data[73][15] <=234;	data[74][15] <=254;	data[75][15] <=240;	data[76][15] <=92;	data[77][15] <=49;	data[78][15] <=85;	data[79][15] <=217;	data[80][15] <=52;	data[81][15] <=239;	data[82][15] <=48;	data[83][15] <=239;	data[84][15] <=178;	data[85][15] <=124;	data[86][15] <=92;	data[87][15] <=97;	data[88][15] <=217;	data[89][15] <=222;	data[90][15] <=103;	data[91][15] <=116;	data[92][15] <=81;	data[93][15] <=211;	data[94][15] <=127;	data[95][15] <=50;	data[96][15] <=38;	data[97][15] <=70;	data[98][15] <=247;	data[99][15] <=156;	data[100][15] <=119;	data[101][15] <=133;	data[102][15] <=256;	data[103][15] <=114;	data[104][15] <=73;	data[105][15] <=31;	data[106][15] <=158;	data[107][15] <=209;	data[108][15] <=55;	data[109][15] <=93;	data[110][15] <=160;	data[111][15] <=163;	data[112][15] <=174;	data[113][15] <=125;	data[114][15] <=229;	data[115][15] <=7;	data[116][15] <=143;	data[117][15] <=91;	data[118][15] <=176;	data[119][15] <=64;	data[120][15] <=193;	data[121][15] <=110;	data[122][15] <=42;	data[123][15] <=180;	data[124][15] <=113;	data[125][15] <=238;	data[126][15] <=144;	data[127][15] <=183;
	
	data[0][0] <=10;	data[1][0] <=38;	data[2][0] <=209;	data[3][0] <=9;
	data[0][1] <=129;	data[1][1] <=38;	data[2][1] <=211;	data[3][1] <=19;
	data[0][2] <=95;	data[1][2] <=2;	data[2][2] <=200;	data[3][2] <=218;
	data[0][3] <=65;	data[1][3] <=18;	data[2][3] <=11;	data[3][3] <=52;
	data[0][4] <=179;	data[1][4] <=207;	data[2][4] <=54;	data[3][4] <=252;
	data[0][5] <=209;	data[1][5] <=74;	data[2][5] <=200;	data[3][5] <=13;
	data[0][6] <=108;	data[1][6] <=167;	data[2][6] <=2;	data[3][6] <=32;
	data[0][7] <=76;	data[1][7] <=41;	data[2][7] <=84;	data[3][7] <=128;
	data[0][8] <=93;	data[1][8] <=42;	data[2][8] <=31;	data[3][8] <=137;
	data[0][9] <=206;	data[1][9] <=180;	data[2][9] <=218;	data[3][9] <=31;
	data[0][10] <=93;	data[1][10] <=114;	data[2][10] <=73;	data[3][10] <=130;
	data[0][11] <=23;	data[1][11] <=8;	data[2][11] <=239;	data[3][11] <=174;
	data[0][12] <=146;	data[1][12] <=195;	data[2][12] <=129;	data[3][12] <=135;
	data[0][13] <=234;	data[1][13] <=252;	data[2][13] <=5;	data[3][13] <=250;
	data[0][14] <=62;	data[1][14] <=177;	data[2][14] <=11;	data[3][14] <=237;
	data[0][15] <=225;	data[1][15] <=70;	data[2][15] <=239;	data[3][15] <=78;
*/

    
    end
    
    
    
    
    
endmodule
